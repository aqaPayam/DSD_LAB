library verilog;
use verilog.vl_types.all;
entity up_down_counter_vlg_vec_tst is
end up_down_counter_vlg_vec_tst;
