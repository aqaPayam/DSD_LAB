library verilog;
use verilog.vl_types.all;
entity pipline_vlg_vec_tst is
end pipline_vlg_vec_tst;
