library verilog;
use verilog.vl_types.all;
entity HW2_vlg_vec_tst is
end HW2_vlg_vec_tst;
